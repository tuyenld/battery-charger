** Profile: "UCC28C42_STEADYSTATE-UCC28C42_SS"  [ e:\sdu-courses\2022-spring\edb2\simulation\ucc28c42_v3\ucc28c42_v3-PSpiceFiles\UCC28C42_STEADYSTATE\UCC28C42_SS.sim ] 

** Creating circuit file "UCC28C42_SS.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../libs/ncp1252.lib" 
.LIB "../../../libs/infineon_simulation model_coolmos_c7_mosfet_650v_spice.lib" 
.LIB "../../../ucc28c42.lib" 
* From [PSPICE NETLIST] section of C:\Users\Dinh-Tuyen Le\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 20m 0m 5ns SKIPBP 
.OPTIONS STEPGMIN
.OPTIONS ABSTOL= 1p
.OPTIONS ITL2= 50
.OPTIONS RELTOL= 0.01
.OPTIONS VNTOL= 1u
.PROBE64 V(*) I(*) D(*) 
.INC "..\UCC28C42_STEADYSTATE.net" 


.END
