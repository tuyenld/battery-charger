** Profile: "UCC28C43_STARTUP-UCC28C43_startup"  [ c:\work\01_ucc28c42\pre-release\01_ucc28c42\02_pspice\modifications after peerreview\ucc28c43_pspice_07nov2008\ucc28c43_pspice_07nov2008\ucc28c43_pspice_trans\ucc28c43-pspicefiles\ucc28c43_startup\ucc28c43_startup.sim ] 

** Creating circuit file "UCC28C43_startup.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../ucc28c43.lib" 
* From [PSPICE NETLIST] section of C:\Cadence\SPB_16.0\tools\PSpice\PSpice.ini file:
.lib "C:\Cadence\SPB_16.0\tools\pspice\library\nom.lib" 

*Analysis directives: 
.TRAN  0 30m 0 {SCHEDULE(0,1000ns,2.5m,25ns)} 
.OPTIONS STEPGMIN
.OPTIONS ABSTOL= 1.0u
.OPTIONS GMIN= 1.0E-11
.OPTIONS ITL4= 10000
.OPTIONS VNTOL= 100.0u
.PROBE V(*) I(*) D(*) 
.INC "..\UCC28C43_STARTUP.net" 


.END
